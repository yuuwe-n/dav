module miniALU(
	input [3:0] op1
	input [3:0] op2
	input operation
	input sign
	); 
	
	
 // The following block contains the logic of your combinational circuit
 always_comb begin
	  // TODO: write the logic for your miniALU here

    end
endmodule 