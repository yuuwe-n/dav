`timescale 1ns/1ns

module miniALU {
    input [3:0] op1;
    input [3:0] op2;
    input [0:0] operation;
    input [0:0] sign;
};

    always_comb

endmodule