`timescale 1ns/1ns

module miniALU_tb ();

	miniALU_top uut(
		.in(send),
		.out(recieve)
	);

endmodule
